module Shift 
#(parameter Width=16)
(
	input  	   [Width-1:0] A,
	input      [2:0] F,
	output reg C,Z,N,P,
	output reg [Width-1:0] Out
);

reg Cshift;

always @(*) 
begin
	case (F)
        3'b000:					//SHL
	    {C,Out} = {A,1'b0};
////////////////////////////////////////////////////////////
        3'b001:					//SHR
	    {Out,C} = {1'b0,A};
////////////////////////////////////////////////////////////
        3'b010:					//SAL
	    {C,Out} = {A,1'b0};
////////////////////////////////////////////////////////////
        3'b011:					//SAR
	    {Out,C} = {A[Width-1],A};
////////////////////////////////////////////////////////////
        3'b100:					//ROL
            {C,Out} = {A,A[Width-1]};
////////////////////////////////////////////////////////////
        3'b101:					//ROR
	    {Out,C} = {A[0],A};
////////////////////////////////////////////////////////////
	3'b110:					//RCL
	begin
	 	Cshift = C;
		{C,Out} = {A,Cshift};
	end      
////////////////////////////////////////////////////////////
	3'b111:					//RCR
	begin
	 	Cshift = C;
		{Out,C} = {Cshift,A};
	end        
////////////////////////////////////////////////////////////                  
        default: 
	begin
            Out = {Width{1'b0}};
            C   = 1'b0;
	    Z 	= 1'b0;
   	    N 	= 1'b0;
    	    P 	= 1'b0;
        end
////////////////////////////////////////////////////////////
        endcase


	Z = ~|Out;		//Zero Flag
    	N = Out[Width-1];	//Negative Flag
    	P = ~^Out;		//Parity Flag
    
end

endmodule
